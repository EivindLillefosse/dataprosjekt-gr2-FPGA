----------------------------------------------------------------------------------
-- Company: NTNU
-- Engineer: Eivind Lillefosse
-- 
-- Create Date: 08.11.2025
-- Design Name: CNN Real Data Testbench
-- Module Name: cnn_real_data_tb - Behavioral
-- Project Name: CNN Accelerator
-- Target Devices: Xilinx FPGA
-- Tool Versions: 
-- Description: Testbench for CNN using real Google Quick Draw or MNIST data
-- 
-- Usage:
--   1. Export test image: python model/export_test_image.py --category apple --index 0
--   2. Run simulation: vivado -mode batch -source scripts/run-single-testbench.tcl -tclargs cnn_real_data
--   3. Compare results: python model/debug_comparison.py --vivado <path> --npz model/intermediate_values.npz
--
-- Dependencies: 
--   - work.test_image_pkg (generated by model/export_test_image.py)
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
use work.types_pkg.all;
use work.test_image_pkg.all;  -- Real test image data from export script

-- Required for file I/O operations
use STD.TEXTIO.ALL;
use IEEE.STD_LOGIC_TEXTIO.ALL;
-- Optional: VHDL-2008 simulator control (std.env). Some simulators support this to stop/finish simulation.
use std.env.all;

entity cnn_real_data_tb is
end cnn_real_data_tb;

architecture Behavioral of cnn_real_data_tb is
    -- Test parameters (matching CNN top-level)
    constant IMAGE_SIZE : integer := 28;
    
    -- Final output will be from CONV_2 with 16 filters
    constant FINAL_NUM_FILTERS : integer := 16;
    
    -- Clock period
    constant CLK_PERIOD : time := 10 ns;
    
    -- UUT signals
    signal clk : STD_LOGIC := '0';
    signal rst : STD_LOGIC := '0';
    
    -- Request/response signals for output
    signal output_req_row   : integer := 0;
    signal output_req_col   : integer := 0;
    signal output_req_valid : std_logic := '0';
    signal output_req_ready : std_logic;
    
    -- Request/response signals for input
    signal input_req_row    : integer;
    signal input_req_col    : integer;
    signal input_req_valid  : std_logic;
    signal input_req_ready  : std_logic := '0';
    
    -- Data signals
    signal input_pixel : WORD_ARRAY_16(0 to 0) := (others => (others => '0'));
    signal input_valid : std_logic := '0';
    signal input_ready : std_logic;
    
    signal output_pixel : WORD_ARRAY_16(0 to FINAL_NUM_FILTERS-1);
    signal output_valid : std_logic;
    signal output_ready : std_logic := '0';
    
    -- DEBUG: Intermediate layer signals
    signal debug_conv1_pixel : WORD_ARRAY_16(0 to 7);  -- 8 filters
    signal debug_conv1_valid : std_logic;
    signal debug_conv1_ready : std_logic := '0';
    signal debug_conv1_row   : natural := 0;
    signal debug_conv1_col   : natural := 0;
    
    signal debug_pool1_pixel : WORD_ARRAY_16(0 to 7);  -- 8 filters
    signal debug_pool1_valid : std_logic;
    signal debug_pool1_ready : std_logic := '0';
    signal debug_pool1_row   : natural := 0;
    signal debug_pool1_col   : natural := 0;
    
    signal debug_conv2_pixel : WORD_ARRAY_16(0 to 15); -- 16 filters
    signal debug_conv2_valid : std_logic;
    signal debug_conv2_ready : std_logic := '0';
    signal debug_conv2_row   : natural := 0;
    signal debug_conv2_col   : natural := 0;
    
    -- Test image data (28x28 image)
    type test_image_type is array (0 to IMAGE_SIZE-1, 0 to IMAGE_SIZE-1) of integer;
    
    -- Function to load real test image from exported package
    function generate_test_image return test_image_type is
        variable temp_image : test_image_type;
    begin
        -- Load real Quick Draw or MNIST data from exported package
        for row in 0 to IMAGE_SIZE-1 loop
            for col in 0 to IMAGE_SIZE-1 loop
                temp_image(row, col) := TEST_IMAGE_DATA(row, col);
            end loop;
        end loop;
        return temp_image;
    end function;
    
    -- Use real test image data
    constant test_image : test_image_type := generate_test_image;
    
    -- Test control signals
    signal test_done : boolean := false;

begin
    -- Unit Under Test (UUT) - CNN Top-Level with debug outputs
    uut: entity work.cnn_top_debug
        generic map (
            IMAGE_SIZE => IMAGE_SIZE
        )
        port map (
            clk              => clk,
            rst              => rst,
            
            -- Output request interface
            output_req_row   => output_req_row,
            output_req_col   => output_req_col,
            output_req_valid => output_req_valid,
            output_req_ready => output_req_ready,
            
            -- Input request interface
            input_req_row    => input_req_row,
            input_req_col    => input_req_col,
            input_req_valid  => input_req_valid,
            input_req_ready  => input_req_ready,
            
            -- Data interfaces
            input_pixel      => input_pixel,
            input_valid      => input_valid,
            input_ready      => input_ready,
            
            output_pixel     => output_pixel,
            output_valid     => output_valid,
            output_ready     => output_ready,
            
            -- DEBUG: Intermediate layer outputs
            debug_conv1_pixel => debug_conv1_pixel,
            debug_conv1_valid => debug_conv1_valid,
            debug_conv1_ready => debug_conv1_ready,
            debug_conv1_row   => debug_conv1_row,
            debug_conv1_col   => debug_conv1_col,
            
            debug_pool1_pixel => debug_pool1_pixel,
            debug_pool1_valid => debug_pool1_valid,
            debug_pool1_ready => debug_pool1_ready,
            debug_pool1_row   => debug_pool1_row,
            debug_pool1_col   => debug_pool1_col,
            
            debug_conv2_pixel => debug_conv2_pixel,
            debug_conv2_valid => debug_conv2_valid,
            debug_conv2_ready => debug_conv2_ready,
            debug_conv2_row   => debug_conv2_row,
            debug_conv2_col   => debug_conv2_col
        );

    -- Clock process
    clk_process: process
    begin
        while not test_done loop
            clk <= '0';
            wait for CLK_PERIOD/2;
            clk <= '1';
            wait for CLK_PERIOD/2;
        end loop;
        wait;
    end process;

    -- Input pixel provider process
    -- Responds to input position requests from the CNN
    input_provider: process(clk)
        variable req_pending : boolean := false;
        variable req_row_buf : integer := 0;
        variable req_col_buf : integer := 0;
    begin
        if rising_edge(clk) then
            if rst = '1' then
                input_req_ready <= '0';
                input_valid <= '0';
                req_pending := false;
            else
                -- Default: not ready for new requests, no data valid
                input_req_ready <= '0';
                input_valid <= '0';
                
                -- Accept new position requests
                if input_req_valid = '1' and not req_pending then
                    input_req_ready <= '1';  -- Acknowledge request
                    req_row_buf := input_req_row;
                    req_col_buf := input_req_col;
                    req_pending := true;
                end if;
                
                -- Provide data for pending request
                if req_pending then
                    if req_row_buf >= 0 and req_row_buf < IMAGE_SIZE and 
                       req_col_buf >= 0 and req_col_buf < IMAGE_SIZE then
                        input_pixel(0) <= std_logic_vector(to_unsigned(test_image(req_row_buf, req_col_buf), 16));
                    else
                        -- Provide zero for out-of-bounds pixels (padding)
                        input_pixel(0) <= (others => '0');
                    end if;
                    input_valid <= '1';
                    
                    -- Wait for acknowledgment
                    if input_ready = '1' then
                        req_pending := false;
                    end if;
                end if;
            end if;
        end if;
    end process;
    
    -- Monitor input requests (separate process for reporting)
    input_monitor: process(clk)
    begin
        if rising_edge(clk) then
            if input_req_valid = '1' and input_req_ready = '1' then
                if input_req_row >= 0 and input_req_row < IMAGE_SIZE and 
                   input_req_col >= 0 and input_req_col < IMAGE_SIZE then
                    report "Input requested [" & integer'image(input_req_row) & "," & integer'image(input_req_col) & "]";
                else
                    report "Input requested (padding) [" & integer'image(input_req_row) & "," & integer'image(input_req_col) & "]";
                end if;
            end if;
            
            if input_valid = '1' and input_ready = '1' then
                report "Input provided: " & integer'image(to_integer(unsigned(input_pixel(0))));
            end if;
        end if;
    end process;

    -- Output monitor process with intermediate value capture
    output_monitor: process(clk)
        file debug_file : text open write_mode is "cnn_intermediate_debug.txt";
        variable debug_line : line;
    begin
        if rising_edge(clk) then
            -- Monitor input requests
            if input_req_valid = '1' and input_req_ready = '1' then
                write(debug_line, string'("INPUT_REQUEST: ["));
                write(debug_line, input_req_row);
                write(debug_line, ',');
                write(debug_line, input_req_col);
                write(debug_line, ']');
                writeline(debug_file, debug_line);
            end if;
            
            -- Monitor input provision
            if input_valid = '1' and input_ready = '1' then
                write(debug_line, string'("INPUT_PROVIDED: ["));
                write(debug_line, input_req_row);  -- Use last requested position
                write(debug_line, ',');
                write(debug_line, input_req_col);
                write(debug_line, string'("] "));
                write(debug_line, to_integer(unsigned(input_pixel(0))));
                writeline(debug_file, debug_line);
            end if;
            
            -- Monitor Conv1 outputs (Layer 0)
            if debug_conv1_valid = '1' then
                write(debug_line, string'("LAYER0_CONV1_OUTPUT: ["));
                write(debug_line, debug_conv1_row);
                write(debug_line, ',');
                write(debug_line, debug_conv1_col);
                write(debug_line, ']');
                writeline(debug_file, debug_line);
                for i in 0 to 7 loop
                    write(debug_line, string'("  Filter_"));
                    write(debug_line, i);
                    write(debug_line, string'(": "));
                    write(debug_line, to_integer(signed(debug_conv1_pixel(i))));
                    writeline(debug_file, debug_line);
                end loop;
                debug_conv1_ready <= '1';
            else
                debug_conv1_ready <= '0';
            end if;
            
            -- Monitor Pool1 outputs (Layer 1)
            if debug_pool1_valid = '1' then
                write(debug_line, string'("LAYER1_POOL1_OUTPUT: ["));
                write(debug_line, debug_pool1_row);
                write(debug_line, ',');
                write(debug_line, debug_pool1_col);
                write(debug_line, ']');
                writeline(debug_file, debug_line);
                for i in 0 to 7 loop
                    write(debug_line, string'("  Filter_"));
                    write(debug_line, i);
                    write(debug_line, string'(": "));
                    write(debug_line, to_integer(signed(debug_pool1_pixel(i))));
                    writeline(debug_file, debug_line);
                end loop;
                debug_pool1_ready <= '1';
            else
                debug_pool1_ready <= '0';
            end if;
            
            -- Monitor Conv2 outputs (Layer 2)
            if debug_conv2_valid = '1' then
                write(debug_line, string'("LAYER2_CONV2_OUTPUT: ["));
                write(debug_line, debug_conv2_row);
                write(debug_line, ',');
                write(debug_line, debug_conv2_col);
                write(debug_line, ']');
                writeline(debug_file, debug_line);
                for i in 0 to 15 loop
                    write(debug_line, string'("  Filter_"));
                    write(debug_line, i);
                    write(debug_line, string'(": "));
                    write(debug_line, to_integer(signed(debug_conv2_pixel(i))));
                    writeline(debug_file, debug_line);
                end loop;
                debug_conv2_ready <= '1';
            else
                debug_conv2_ready <= '0';
            end if;
            
            -- Monitor final outputs (Layer 3 - Pool2)
            if output_valid = '1' and output_ready = '1' then
                report "CNN Output received";
                
                -- CNN_OUTPUT header
                write(debug_line, string'("CNN_OUTPUT: ["));
                write(debug_line, output_req_row);  -- Use requested output position
                write(debug_line, ',');
                write(debug_line, output_req_col);
                write(debug_line, ']');
                writeline(debug_file, debug_line);
                
                for i in 0 to FINAL_NUM_FILTERS-1 loop
                    report "  Filter " & integer'image(i) & ": " & 
                        integer'image(to_integer(signed(output_pixel(i))));
                    -- Write filter output
                    write(debug_line, string'("  Filter_"));
                    write(debug_line, i);
                    write(debug_line, string'(": "));
                    write(debug_line, to_integer(signed(output_pixel(i))));
                    writeline(debug_file, debug_line);
                end loop;
            end if;
        end if;
    end process;

    -- Main test process
    test_process: process
        constant FINAL_OUTPUT_SIZE : integer := 5;  -- After Conv1(26x26)->Pool1(13x13)->Conv2(11x11)->Pool2(5x5)
    begin
        -- Initialize
        rst <= '1';
        output_req_valid <= '0';
        output_ready <= '0';
        
        wait for CLK_PERIOD * 2;
        rst <= '0';
        
        wait for CLK_PERIOD * 2;
        
        report "========================================";
        report "CNN Real Data Test - Starting";
        report "========================================";
        report "Test Image Category: " & TEST_IMAGE_CATEGORY;
        report "Expected Label: " & integer'image(TEST_IMAGE_LABEL);
        report "Image Size: " & integer'image(TEST_IMAGE_SIZE) & "x" & integer'image(TEST_IMAGE_SIZE);
        report "========================================";
        
        report "Test image loaded - sample pixel values:";
        report "  [0,0]=" & integer'image(test_image(0,0)) & 
               "  [0,13]=" & integer'image(test_image(0,13)) & 
               "  [0,27]=" & integer'image(test_image(0,27));
        report "  [13,0]=" & integer'image(test_image(13,0)) & 
               "  [13,13]=" & integer'image(test_image(13,13)) & 
               "  [13,27]=" & integer'image(test_image(13,27));
        report "  [27,0]=" & integer'image(test_image(27,0)) & 
               "  [27,13]=" & integer'image(test_image(27,13)) & 
               "  [27,27]=" & integer'image(test_image(27,27));
        
        -- Request all output positions (5x5 final output)
        for out_row in 0 to FINAL_OUTPUT_SIZE-1 loop
            for out_col in 0 to FINAL_OUTPUT_SIZE-1 loop
                report "Requesting CNN output position [" & integer'image(out_row) & "," & integer'image(out_col) & "]";
                
                -- Send output position request (robust handshake)
                output_req_row <= out_row;
                output_req_col <= out_col;
                output_req_valid <= '1';

                -- Let DUT sample the valid (wait one clock edge)
                wait until rising_edge(clk);

                -- Wait until DUT asserts ready (may be pulsed after sampling)
                while output_req_ready /= '1' loop
                    wait until rising_edge(clk);
                end loop;

                -- Clear request on next clock edge (single-cycle pulse)
                wait until rising_edge(clk);
                output_req_valid <= '0';
                
                -- Wait for output to be ready, then accept it
                -- Set ready high BEFORE the clock edge where output_valid is '1'
                loop
                    -- Pre-assert output_ready
                    output_ready <= '1';
                    wait until rising_edge(clk);
                    -- Check if output was valid on this edge
                    if output_valid = '1' then
                        exit;  -- Both signals were high, monitor will capture
                    end if;
                end loop;
                
                -- Clear ready on next cycle
                output_ready <= '0';
                
                -- Small gap before next request
                wait for CLK_PERIOD;
            end loop;
        end loop;
        
        report "========================================";
        report "All CNN outputs received!";
        report "Category: " & TEST_IMAGE_CATEGORY & " (label " & integer'image(TEST_IMAGE_LABEL) & ")";
        report "========================================";
        
        -- Wait a few more cycles
        wait for CLK_PERIOD * 10;
        
        -- Test reset functionality
        report "Testing CNN reset functionality...";
        rst <= '1';
        wait for CLK_PERIOD * 2;
        rst <= '0';
        
        wait for CLK_PERIOD * 5;
        
        -- Test second run (just first output position)
        report "Testing second CNN run (first position only)...";
        
        output_req_row <= 0;
        output_req_col <= 0;
        output_req_valid <= '1';

        -- Give DUT a clock to sample the request
        wait until rising_edge(clk);

        -- Wait for acknowledgement
        while output_req_ready /= '1' loop
            wait until rising_edge(clk);
        end loop;

        wait until rising_edge(clk);
        output_req_valid <= '0';
        
        -- Fixed handshake for second run too (same pattern)
        loop
            output_ready <= '1';
            wait until rising_edge(clk);
            if output_valid = '1' then
                exit;
            end if;
        end loop;
        output_ready <= '0';
        
        report "Second CNN run completed!";
        
        wait for CLK_PERIOD * 10;
        
        test_done <= true;
        report "========================================";
        report " CNN Real Data Test PASSED";
        report "Category: " & TEST_IMAGE_CATEGORY;
        report "Expected Label: " & integer'image(TEST_IMAGE_LABEL);
        report "========================================";
        
        -- Allow signals to settle for one clock period
        wait for CLK_PERIOD;
        -- Explicitly stop simulation when the simulator supports VHDL-2008 std.env
        -- This forces immediate termination; remove/comment out if your simulator doesn't support std.env
        std.env.stop(0);
        wait;
    end process;

    -- Timeout watchdog
    timeout_watchdog: process
    begin
        -- Simple watchdog pattern used by other testbenches in this repo
        wait for 2000 ms;  -- Longer timeout for full CNN
        if not test_done then
            report "CNN REAL DATA TEST TIMEOUT - Test did not complete within expected time" severity failure;
        end if;
        wait;
    end process;

end Behavioral;
