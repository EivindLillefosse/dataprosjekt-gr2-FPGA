----------------------------------------------------------------------------------
-- Company: NTNU
-- Engineer: 
-- 
-- Create Date: 11.04.2025
-- Design Name: Fully Connected Layer
-- Module Name: Calc Index
-- Project Name: CNN Accelerator
-- Description:  Calculate flattened index from 3D tensor indices
-- 
----------------------------------------------------------------------------------

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
use work.types_pkg.all;
use work.bias_pkg.all;

entity calc_index is
    generic (
        NODES_IN       : integer := 400;
        INPUT_CHANNELS : integer := 16;
        INPUT_SIZE     : integer := 5
    );
    port (
        clk     : in  std_logic;
        rst     : in  std_logic;
        enable  : in  std_logic;  -- Start requesting pixels
        
        -- Request to upstream (max pooling layer) - only row/col needed
        req_row     : out integer; -- plain integer to match top-level signals
        req_col     : out integer; -- plain integer to match top-level signals
        req_valid   : out std_logic;
        
        -- Input from max pooling: all 16 channels at once (16x8 bits)
        pool_pixel_data  : in WORD_ARRAY_16(0 to INPUT_CHANNELS-1);
        pool_pixel_valid : in std_logic;
        pool_pixel_ready : out std_logic;
        
        -- Output to FC layer: selected single channel pixel
        fc_pixel_out    : out WORD_16;
        fc_pixel_valid  : out std_logic;
        fc_pixel_ready  : in  std_logic;
        
        -- Current index being requested (for debugging/monitoring)
        curr_index  : out integer range 0 to NODES_IN-1;
        
        -- Done signal when all 400 pixels requested
        done        : out std_logic
    );
end calc_index;

architecture Structural of calc_index is
    constant NUM_POSITIONS                         : integer := INPUT_SIZE * INPUT_SIZE;  -- 25 spatial positions
    
    signal position_counter                        : integer range 0 to NUM_POSITIONS-1 := 0;
    attribute keep_pos_cnt                         : string;
    attribute keep_pos_cnt of position_counter     : signal is "true";
    attribute syn_keep_pos_cnt                     : string;
    attribute syn_keep_pos_cnt of position_counter : signal is "true";
    signal channel_counter                         : integer range 0 to INPUT_CHANNELS-1 := 0;
    attribute keep_chan_cnt                        : string;
    attribute keep_chan_cnt of channel_counter     : signal is "true";
    attribute syn_keep_chan_cnt                    : string;
    attribute syn_keep_chan_cnt of channel_counter : signal is "true";
    signal internal_done                           : std_logic := '0';
    signal pool_data_captured                      : WORD_ARRAY_16(0 to INPUT_CHANNELS-1) := (others => (others => '0'));
    signal data_valid                              : std_logic := '0';
    signal last_chan                               : std_logic := '0';
    -- Registered outputs for request coordinates to preserve in synthesis
    signal req_row_reg : integer                   := 0;
    attribute keep_req_row_reg                     : string;
    attribute keep_req_row_reg of req_row_reg      : signal is "true";
    attribute syn_keep_req_row_reg                 : string;
    attribute syn_keep_req_row_reg of req_row_reg  : signal is "true";
    signal req_col_reg : integer                   := 0;
    attribute keep_req_col_reg                     : string;
    attribute keep_req_col_reg of req_col_reg      : signal is "true";
    attribute syn_keep_req_col_reg                 : string;
    attribute syn_keep_req_col_reg of req_col_reg  : signal is "true";
begin
    
    -- Main state machine: request Pool2 position, capture 16 channels, send to FC1 sequentially
    process(clk)
    begin
        if rising_edge(clk) then
            if rst = '1' then
                position_counter <= 0;
                channel_counter   <= 0;
                internal_done    <= '0';
                data_valid       <= '0';
                pool_data_captured <= (others => (others => '0'));
                last_chan        <= '0';
                req_row_reg      <= 0;
                req_col_reg      <= 0;
            elsif enable = '1' then
                if internal_done = '1' then
                    -- Restart
                    position_counter   <= 0;
                    channel_counter    <= 0;
                    internal_done      <= '0';
                    data_valid         <= '0';
                    pool_data_captured <= (others => (others => '0'));
                    last_chan          <= '0';
                    req_row_reg        <= 0;
                    req_col_reg        <= 0;
                else
                    -- When Pool2 delivers data, capture it and start sending channels
                    if pool_pixel_valid = '1' and data_valid = '0' then
                        pool_data_captured <= pool_pixel_data;
                        data_valid         <= '1';
                        channel_counter    <= 0;
                    end if;
                    
                    if channel_counter = INPUT_CHANNELS - 1 then 
                        last_chan <= '1';
                    end if;
                    
                    -- Send captured channels sequentially to FC1
                    if data_valid = '1' and fc_pixel_ready = '1' then

                        if channel_counter < INPUT_CHANNELS - 1 then
                            -- Move to next channel
                            channel_counter <= channel_counter + 1;
                        else
                            -- Sent all 16 channels for this position
                            channel_counter <= 0;
                            data_valid <= '0';
                            last_chan <= '0';
                            
                            if position_counter = NUM_POSITIONS - 1 then
                                -- All positions done (we just finished the last position)
                                internal_done <= '1';
                            else
                                -- Move to next position and update row/col incrementally
                                position_counter <= position_counter + 1;
                                if req_col_reg = INPUT_SIZE - 1 then
                                    req_col_reg <= 0;
                                    req_row_reg <= req_row_reg + 1;
                                else
                                    req_col_reg <= req_col_reg + 1;
                                end if;
                            end if;
                        end if;
                    elsif position_counter = NUM_POSITIONS - 1 and last_chan = '1' then
                        internal_done <= '1';
                    end if;
                end if;
            elsif enable = '0' then
                internal_done <= '0';
                data_valid    <= '0';
            end if;
        end if;
    end process;
    
    -- Reverse calculation: position to 2D coordinates
    -- position = row * INPUT_SIZE + col
    req_row     <= req_row_reg;
    req_col     <= req_col_reg;
    req_valid   <= enable and not internal_done and not data_valid;  -- Only request when not processing channels

    -- Output current channel from captured data
    fc_pixel_out   <= pool_data_captured(channel_counter);
    fc_pixel_valid <= data_valid and enable and not internal_done;
    
    -- Assert ready when waiting for Pool2 data
    pool_pixel_ready <= enable and not internal_done and not data_valid;
    
    -- Status outputs
    curr_index  <= position_counter * INPUT_CHANNELS + channel_counter;  -- Absolute pixel index (0-399)
    done        <= internal_done;

end architecture Structural;