library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

package bias_pkg is
    type layer_0_conv2d_t is array(0 to 29) of signed(7 downto 0);
    constant layer_0_conv2d_BIAS : layer_0_conv2d_t := (
        0 => to_signed(-1, 8),
        1 => to_signed(-8, 8),
        2 => to_signed(-19, 8),
        3 => to_signed(4, 8),
        4 => to_signed(-4, 8),
        5 => to_signed(-8, 8),
        6 => to_signed(0, 8),
        7 => to_signed(-8, 8),
        8 => to_signed(-12, 8),
        9 => to_signed(-3, 8),
        10 => to_signed(-13, 8),
        11 => to_signed(-4, 8),
        12 => to_signed(11, 8),
        13 => to_signed(-2, 8),
        14 => to_signed(-1, 8),
        15 => to_signed(-15, 8),
        16 => to_signed(-18, 8),
        17 => to_signed(-11, 8),
        18 => to_signed(-21, 8),
        19 => to_signed(-1, 8),
        20 => to_signed(-1, 8),
        21 => to_signed(-8, 8),
        22 => to_signed(-10, 8),
        23 => to_signed(-7, 8),
        24 => to_signed(-1, 8),
        25 => to_signed(-14, 8),
        26 => to_signed(5, 8),
        27 => to_signed(2, 8),
        28 => to_signed(3, 8),
        29 => to_signed(0, 8)
    );
    type layer_2_conv2d_1_t is array(0 to 59) of signed(7 downto 0);
    constant layer_2_conv2d_1_BIAS : layer_2_conv2d_1_t := (
        0 => to_signed(-2, 8),
        1 => to_signed(-5, 8),
        2 => to_signed(-2, 8),
        3 => to_signed(-10, 8),
        4 => to_signed(1, 8),
        5 => to_signed(6, 8),
        6 => to_signed(-6, 8),
        7 => to_signed(-7, 8),
        8 => to_signed(-1, 8),
        9 => to_signed(-4, 8),
        10 => to_signed(3, 8),
        11 => to_signed(-2, 8),
        12 => to_signed(-1, 8),
        13 => to_signed(-7, 8),
        14 => to_signed(-5, 8),
        15 => to_signed(1, 8),
        16 => to_signed(-8, 8),
        17 => to_signed(-3, 8),
        18 => to_signed(-3, 8),
        19 => to_signed(1, 8),
        20 => to_signed(-4, 8),
        21 => to_signed(0, 8),
        22 => to_signed(-2, 8),
        23 => to_signed(-11, 8),
        24 => to_signed(-1, 8),
        25 => to_signed(-8, 8),
        26 => to_signed(4, 8),
        27 => to_signed(-12, 8),
        28 => to_signed(5, 8),
        29 => to_signed(-1, 8),
        30 => to_signed(-11, 8),
        31 => to_signed(-7, 8),
        32 => to_signed(-2, 8),
        33 => to_signed(-10, 8),
        34 => to_signed(-10, 8),
        35 => to_signed(-2, 8),
        36 => to_signed(-6, 8),
        37 => to_signed(-5, 8),
        38 => to_signed(-2, 8),
        39 => to_signed(-5, 8),
        40 => to_signed(-4, 8),
        41 => to_signed(-6, 8),
        42 => to_signed(-2, 8),
        43 => to_signed(-10, 8),
        44 => to_signed(-13, 8),
        45 => to_signed(-1, 8),
        46 => to_signed(-12, 8),
        47 => to_signed(-4, 8),
        48 => to_signed(-2, 8),
        49 => to_signed(-1, 8),
        50 => to_signed(-1, 8),
        51 => to_signed(-2, 8),
        52 => to_signed(-4, 8),
        53 => to_signed(-5, 8),
        54 => to_signed(-12, 8),
        55 => to_signed(-2, 8),
        56 => to_signed(8, 8),
        57 => to_signed(-1, 8),
        58 => to_signed(-4, 8),
        59 => to_signed(-2, 8)
    );
    type layer_5_dense_t is array(0 to 119) of signed(7 downto 0);
    constant layer_5_dense_BIAS : layer_5_dense_t := (
        0 => to_signed(-2, 8),
        1 => to_signed(0, 8),
        2 => to_signed(-4, 8),
        3 => to_signed(-1, 8),
        4 => to_signed(-2, 8),
        5 => to_signed(-2, 8),
        6 => to_signed(0, 8),
        7 => to_signed(-3, 8),
        8 => to_signed(-1, 8),
        9 => to_signed(-1, 8),
        10 => to_signed(-2, 8),
        11 => to_signed(-3, 8),
        12 => to_signed(-2, 8),
        13 => to_signed(0, 8),
        14 => to_signed(-2, 8),
        15 => to_signed(0, 8),
        16 => to_signed(-3, 8),
        17 => to_signed(-2, 8),
        18 => to_signed(-1, 8),
        19 => to_signed(-1, 8),
        20 => to_signed(-3, 8),
        21 => to_signed(5, 8),
        22 => to_signed(-3, 8),
        23 => to_signed(-1, 8),
        24 => to_signed(-1, 8),
        25 => to_signed(-2, 8),
        26 => to_signed(-1, 8),
        27 => to_signed(0, 8),
        28 => to_signed(-4, 8),
        29 => to_signed(-2, 8),
        30 => to_signed(-3, 8),
        31 => to_signed(1, 8),
        32 => to_signed(-3, 8),
        33 => to_signed(-1, 8),
        34 => to_signed(-1, 8),
        35 => to_signed(-1, 8),
        36 => to_signed(-2, 8),
        37 => to_signed(1, 8),
        38 => to_signed(2, 8),
        39 => to_signed(-1, 8),
        40 => to_signed(-1, 8),
        41 => to_signed(-1, 8),
        42 => to_signed(-1, 8),
        43 => to_signed(-5, 8),
        44 => to_signed(0, 8),
        45 => to_signed(-3, 8),
        46 => to_signed(-3, 8),
        47 => to_signed(-2, 8),
        48 => to_signed(0, 8),
        49 => to_signed(-2, 8),
        50 => to_signed(-2, 8),
        51 => to_signed(-2, 8),
        52 => to_signed(-4, 8),
        53 => to_signed(-5, 8),
        54 => to_signed(-2, 8),
        55 => to_signed(2, 8),
        56 => to_signed(1, 8),
        57 => to_signed(-5, 8),
        58 => to_signed(4, 8),
        59 => to_signed(-2, 8),
        60 => to_signed(2, 8),
        61 => to_signed(-1, 8),
        62 => to_signed(-4, 8),
        63 => to_signed(-2, 8),
        64 => to_signed(1, 8),
        65 => to_signed(-3, 8),
        66 => to_signed(-1, 8),
        67 => to_signed(-4, 8),
        68 => to_signed(-3, 8),
        69 => to_signed(-4, 8),
        70 => to_signed(-3, 8),
        71 => to_signed(-2, 8),
        72 => to_signed(3, 8),
        73 => to_signed(-4, 8),
        74 => to_signed(-2, 8),
        75 => to_signed(-4, 8),
        76 => to_signed(-1, 8),
        77 => to_signed(-3, 8),
        78 => to_signed(2, 8),
        79 => to_signed(-2, 8),
        80 => to_signed(6, 8),
        81 => to_signed(-2, 8),
        82 => to_signed(-1, 8),
        83 => to_signed(-2, 8),
        84 => to_signed(-2, 8),
        85 => to_signed(2, 8),
        86 => to_signed(0, 8),
        87 => to_signed(-1, 8),
        88 => to_signed(-1, 8),
        89 => to_signed(-1, 8),
        90 => to_signed(4, 8),
        91 => to_signed(-3, 8),
        92 => to_signed(-3, 8),
        93 => to_signed(-3, 8),
        94 => to_signed(-2, 8),
        95 => to_signed(-4, 8),
        96 => to_signed(-2, 8),
        97 => to_signed(2, 8),
        98 => to_signed(-1, 8),
        99 => to_signed(-1, 8),
        100 => to_signed(5, 8),
        101 => to_signed(-4, 8),
        102 => to_signed(-1, 8),
        103 => to_signed(-2, 8),
        104 => to_signed(-1, 8),
        105 => to_signed(-2, 8),
        106 => to_signed(1, 8),
        107 => to_signed(-1, 8),
        108 => to_signed(-2, 8),
        109 => to_signed(-4, 8),
        110 => to_signed(2, 8),
        111 => to_signed(-4, 8),
        112 => to_signed(-3, 8),
        113 => to_signed(-3, 8),
        114 => to_signed(2, 8),
        115 => to_signed(6, 8),
        116 => to_signed(3, 8),
        117 => to_signed(-3, 8),
        118 => to_signed(0, 8),
        119 => to_signed(-2, 8)
    );
    type layer_6_dense_1_t is array(0 to 19) of signed(7 downto 0);
    constant layer_6_dense_1_BIAS : layer_6_dense_1_t := (
        0 => to_signed(11, 8),
        1 => to_signed(-5, 8),
        2 => to_signed(6, 8),
        3 => to_signed(10, 8),
        4 => to_signed(-5, 8),
        5 => to_signed(-3, 8),
        6 => to_signed(-2, 8),
        7 => to_signed(0, 8),
        8 => to_signed(-6, 8),
        9 => to_signed(6, 8),
        10 => to_signed(-4, 8),
        11 => to_signed(-8, 8),
        12 => to_signed(2, 8),
        13 => to_signed(7, 8),
        14 => to_signed(1, 8),
        15 => to_signed(-3, 8),
        16 => to_signed(-5, 8),
        17 => to_signed(-6, 8),
        18 => to_signed(6, 8),
        19 => to_signed(-5, 8)
    );
end package bias_pkg;

package body bias_pkg is
end package body bias_pkg;
