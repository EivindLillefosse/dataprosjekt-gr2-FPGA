-- Test vectors for convolution debugging
-- Simple 3x3 pattern for verification

constant test_pattern : test_image_type := (
    (1, 2, 3),
    (4, 5, 6),
    (7, 8, 9)
);
